// Created by prof. Mingu Kang @VVIP Lab in UCSD ECE department
// Modified for ECE284 Part B Requirements
`timescale 1ns/1ps

module core_tb;

parameter bw       = 4;
parameter psum_bw  = 16;
parameter len_kij  = 9;
parameter len_onij = 4; 
parameter col      = 8;
parameter row      = 8;
parameter len_nij  = 4;

reg clk   = 0;
reg reset = 1;

wire [33:0] inst_q;

reg [bw*row-1:0] D_xmem_q = 0;

// XMEM control
reg CEN_xmem = 1;
reg WEN_xmem = 1;
reg [10:0] A_xmem = 0;
reg CEN_xmem_q = 1;
reg WEN_xmem_q = 1;
reg [10:0] A_xmem_q = 0;

// PMEM control
reg CEN_pmem = 1;
reg WEN_pmem = 1;
reg [10:0] A_pmem = 0;
reg CEN_pmem_q = 1;
reg WEN_pmem_q = 1;
reg [10:0] A_pmem_q = 0;

// control to FIFOs / core
reg ofifo_rd_q = 0;
reg ififo_wr_q = 0;
reg ififo_rd_q = 0;
reg l0_rd_q    = 0;
reg l0_wr_q    = 0;
reg execute_q  = 0;
reg load_q     = 0;
reg acc_q      = 0;
reg acc        = 0;

// unregistered drivers
reg [bw*row-1:0] D_xmem;
reg [psum_bw*col-1:0] answer;

reg ofifo_rd;
reg ififo_wr;
reg ififo_rd;
reg l0_rd;
reg l0_wr;
reg execute;
reg load;

wire ofifo_valid;
wire [col*psum_bw-1:0] sfp_out;

// file handles
integer x_file, x_scan_file;
integer w_file, w_scan_file;
integer acc_file, acc_scan_file;
integer out_file, out_scan_file;
integer captured_data;
integer t, i, j, kij;
integer error;

// pack instruction bus
assign inst_q[33]    = acc_q;
assign inst_q[32]    = CEN_pmem_q;
assign inst_q[31]    = WEN_pmem_q;
assign inst_q[30:20] = A_pmem_q;
assign inst_q[19]    = CEN_xmem_q;
assign inst_q[18]    = WEN_xmem_q;
assign inst_q[17:7]  = A_xmem_q;
assign inst_q[6]     = ofifo_rd_q;
assign inst_q[5]     = ififo_wr_q;
assign inst_q[4]     = ififo_rd_q;
assign inst_q[3]     = l0_rd_q;
assign inst_q[2]     = l0_wr_q;
assign inst_q[1]     = execute_q;
assign inst_q[0]     = load_q;

// ---------------------------------------------
// core instance
// ---------------------------------------------
core #(
  .bw(bw),
  .col(col),
  .row(row)
) core_instance (
  .clk     (clk),
  .inst    (inst_q),
  .ofifo_valid(ofifo_valid),
  .D_xmem  (D_xmem_q),
  .sfp_out (sfp_out),
  .reset   (reset),
  .mode    (1'b0) 
);

// ---------------------------------------------
// main test sequence
// ---------------------------------------------
initial begin
  $dumpfile("core_tb.vcd");
  $dumpvars(0, core_tb);

  // initialize default values
  D_xmem   = 0;
  CEN_xmem = 1;
  WEN_xmem = 1;
  A_xmem   = 0;

  A_pmem   = 0;
  CEN_pmem = 1;
  WEN_pmem = 1;

  ofifo_rd = 0;
  ififo_wr = 0;
  ififo_rd = 0;
  l0_rd    = 0;
  l0_wr    = 0;
  execute  = 0;
  load     = 0;
  acc      = 0;

  // -------------------------
  // system reset
  // -------------------------
  #0.5 clk = 1'b0; reset = 1;
  #0.5 clk = 1'b1;

  for (i=0; i<10; i=i+1) begin
    #0.5 clk = 1'b0;
    #0.5 clk = 1'b1;
  end

  #0.5 clk = 1'b0; reset = 0;
  #0.5 clk = 1'b1;

  #0.5 clk = 1'b0;
  #0.5 clk = 1'b1;

  // -------------------------
  // load activation into XMEM

  x_file = $fopen("input.txt", "r"); 
  x_scan_file = $fscanf(x_file,"%s", captured_data);
  x_scan_file = $fscanf(x_file,"%s", captured_data);
  x_scan_file = $fscanf(x_file,"%s", captured_data);

  for (t=0; t<len_nij; t=t+1) begin
    #0.5 clk = 1'b0;
      x_scan_file = $fscanf(x_file,"%32b", D_xmem);
      WEN_xmem = 0;
      CEN_xmem = 0;
      if (t>0) A_xmem = A_xmem + 1;
    #0.5 clk = 1'b1;
  end

  #0.5 clk = 1'b0;
    WEN_xmem = 1;
    CEN_xmem = 1;
    A_xmem   = 0;
  #0.5 clk = 1'b1;

  $fclose(x_file);

  w_file = $fopen("weight.txt", "r");
  w_scan_file = $fscanf(w_file,"%s", captured_data);
  w_scan_file = $fscanf(w_file,"%s", captured_data);
  w_scan_file = $fscanf(w_file,"%s", captured_data);

  // -------------------------
  // kij loop (3x3 kernel)
  // -------------------------
  A_pmem = 0; // pmem write pointer for partial sums

  for (kij=0; kij<len_kij; kij=kij+1) begin

    // kernel loop reset
    #0.5 clk = 1'b0; reset = 1;
    #0.5 clk = 1'b1;

    for (i=0; i<10; i=i+1) begin
      #0.5 clk = 1'b0;
      #0.5 clk = 1'b1;
    end

    #0.5 clk = 1'b0; reset = 0;
    #0.5 clk = 1'b1;

    #0.5 clk = 1'b0;
    #0.5 clk = 1'b1;

    // -------------------------
    // write kernel weights to XMEM
    // base address for kernel
    // -------------------------
    A_xmem = 11'b10000000000;

    for (t=0; t<col; t=t+1) begin
      #0.5 clk = 1'b0;
        w_scan_file = $fscanf(w_file,"%32b", D_xmem);
        WEN_xmem = 0;
        CEN_xmem = 0;
        if (t>0) A_xmem = A_xmem + 1;
      #0.5 clk = 1'b1;
    end

    #0.5 clk = 1'b0;
      WEN_xmem = 1;
      CEN_xmem = 1;
      A_xmem   = 0;
    #0.5 clk = 1'b1;

    // -------------------------
    // kernel data XMEM -> L0
    // -------------------------
    A_xmem = 11'b10000000000;
    for (t=0; t<col; t=t+1) begin
      #0.5 clk = 1'b0;
        CEN_xmem = 0;
        WEN_xmem = 1;
        l0_wr    = 1;
        if (t>0) A_xmem = A_xmem + 1;
      #0.5 clk = 1'b1;
    end

    #0.5 clk = 1'b0;
      CEN_xmem = 1;
      l0_wr    = 0;
    #0.5 clk = 1'b1;

    // -------------------------
    // kernel loading to PEs
    // -------------------------
    for (t=0; t<col; t=t+1) begin
      #0.5 clk = 1'b0;
        l0_rd = 1;
        load  = 1;
      #0.5 clk = 1'b1;
    end

    #0.5 clk = 1'b0;
      l0_rd = 0;
      load  = 0;
    #0.5 clk = 1'b1;

    // -------------------------
    // intermission
    // -------------------------
    #0.5 clk = 1'b0;
      load  = 0;
      l0_rd = 0;
    #0.5 clk = 1'b1;

    for (i=0; i<10; i=i+1) begin
      #0.5 clk = 1'b0;
      #0.5 clk = 1'b1;
    end

    // -------------------------
    // activation XMEM -> L0
    // -------------------------
    A_xmem = 0;
    for (t=0; t<len_nij; t=t+1) begin
      #0.5 clk = 1'b0;
        CEN_xmem = 0;
        WEN_xmem = 1;
        l0_wr    = 1;
        if (t>0) A_xmem = A_xmem + 1;
      #0.5 clk = 1'b1;
    end

    #0.5 clk = 1'b0;
      CEN_xmem = 1;
      l0_wr    = 0;
    #0.5 clk = 1'b1;

    // -------------------------
    // execution
    // -------------------------
    for (t=0; t<len_nij; t=t+1) begin
      #0.5 clk = 1'b0;
        l0_rd    = 1;
        execute = 1;
      #0.5 clk = 1'b1;
    end

    #0.5 clk = 1'b0;
      l0_rd    = 0;
      execute = 0;
    #0.5 clk = 1'b1;

    // -------------------------
    // OFIFO read -> PMEM write
    // -------------------------
    for (t=0; t<len_onij; t=t+1) begin
      #0.5 clk = 1'b0;
        ofifo_rd = 1;
        CEN_pmem = 0;
        WEN_pmem = 0;
      #0.5 clk = 1'b1;
      A_pmem = A_pmem + 1;
    end

    #0.5 clk = 1'b0;
      ofifo_rd = 0;
      CEN_pmem = 1;
      WEN_pmem = 1;
    #0.5 clk = 1'b1;

  end // end of kij loop

  $fclose(w_file); // 

  // -------------------------
  // accumulation & verification
  // -------------------------
  out_file = $fopen("output.txt", "r"); 
  out_scan_file = $fscanf(out_file,"%s", answer);
  out_scan_file = $fscanf(out_file,"%s", answer);
  out_scan_file = $fscanf(out_file,"%s", answer);

  error    = 0;
  acc_file = $fopen("acc_address.txt", "r");

  $display("############ Verification Start #############");

  for (i=0; i<len_onij+1; i=i+1) begin

    #0.5 clk = 1'b0;
    #0.5 clk = 1'b1;

    if (i>0) begin
      out_scan_file = $fscanf(out_file,"%128b", answer);
      if (sfp_out == answer) begin
        $display("%2d-th output featuremap Data matched! :D", i);
      end else begin
        $display("%2d-th output featuremap Data ERROR!!", i);
        $display("sfpout: %128b", sfp_out);
        $display("answer: %128b", answer);
        error = 1;
      end
    end

    // accumulation phase for next output
    #0.5 clk = 1'b0; reset = 1;
    #0.5 clk = 1'b1;
    #0.5 clk = 1'b0; reset = 0;
    #0.5 clk = 1'b1;

    for (j=0; j<len_kij+1; j=j+1) begin
      #0.5 clk = 1'b0;
        if (j < len_kij) begin
          CEN_pmem = 0;
          WEN_pmem = 1;
          acc_scan_file = $fscanf(acc_file,"%11b", A_pmem);
        end else begin
          CEN_pmem = 1;
          WEN_pmem = 1;
        end

        if (j > 0) acc = 1;
      #0.5 clk = 1'b1;
    end

    #0.5 clk = 1'b0; acc = 0;
    #0.5 clk = 1'b1;
  end

  if (error == 0) begin
    $display("############ No error detected ##############");
  end else begin
    $display("############ ERRORS DETECTED ##############");
  end

  $fclose(out_file);
  $fclose(acc_file);

  #10 $finish;

end

always @ (posedge clk) begin
   D_xmem_q   <= D_xmem;
   CEN_xmem_q <= CEN_xmem;
   WEN_xmem_q <= WEN_xmem;
   A_pmem_q   <= A_pmem;
   CEN_pmem_q <= CEN_pmem;
   WEN_pmem_q <= WEN_pmem;
   A_xmem_q   <= A_xmem;
   ofifo_rd_q <= ofifo_rd;
   acc_q      <= acc;
   ififo_wr_q <= ififo_wr;
   ififo_rd_q <= ififo_rd;
   l0_rd_q    <= l0_rd;
   l0_wr_q    <= l0_wr ;
   execute_q  <= execute;
   load_q     <= load;
end

endmodule